module fifo_async #(
    parameters
) (
    port_list
);
    
endmodule