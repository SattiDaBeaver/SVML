module spi_slave #(
    parameter WIDTH = 8;
) (
    input  logic    sclk;
);
    
endmodule